`timescale 1ns / 1ps

//Basic 32 bit decoder, used for instruction input to get registers 
module reg_decoder(
    input [4:0] in,
    output reg [31:0] out
    );
    
    always @ (in) begin
        case(in)
            5'b00000: out = 32'h00000001;
            5'b00001: out = 32'h00000002;
            5'b00010: out = 32'h00000004;
            5'b00011: out = 32'h00000008;
            5'b00100: out = 32'h00000010;
            5'b00101: out = 32'h00000020;
            5'b00110: out = 32'h00000040;
            5'b00111: out = 32'h00000080;
            5'b01000: out = 32'h00000100;
            5'b01001: out = 32'h00000200;
            5'b01010: out = 32'h00000400;
            5'b01011: out = 32'h00000800;
            5'b01100: out = 32'h00001000;
            5'b01101: out = 32'h00002000; 
            5'b01110: out = 32'h00004000;
            5'b01111: out = 32'h00008000;
            5'b10000: out = 32'h00010000;
            5'b10001: out = 32'h00020000;
            5'b10010: out = 32'h00040000;
            5'b10011: out = 32'h00080000;
            5'b10100: out = 32'h00100000;
            5'b10101: out = 32'h00200000;
            5'b10110: out = 32'h00400000;
            5'b10111: out = 32'h00800000;
            5'b11000: out = 32'h01000000;
            5'b11001: out = 32'h02000000;
            5'b11010: out = 32'h04000000;
            5'b11011: out = 32'h08000000;
            5'b11100: out = 32'h10000000;
            5'b11101: out = 32'h20000000;
            5'b11110: out = 32'h40000000;
            5'b11111: out = 32'h80000000;
        endcase
    end
endmodule
