`timescale 1ns / 1ps

//ALU, named Lab 1 because I didn't know we were reusing lab code back then 
//Partially taken from sample code by Northeastern University 
module Lab1 (d, Cout, V, a, b, Cin, S, Z);
   output[31:0] d;
   output Cout, V;
   output reg Z;
   input [31:0] a, b;
   input Cin;
   input [2:0] S;
   
   wire [31:0] c, g, p;
   wire gout, pout;
   
   alu_cell mycell[31:0] (
      .d(d),
      .g(g),
      .p(p),
      .a(a),
      .b(b),
      .c(c),
      .S(S)
   );
   
   lac5 lac(
      .c(c),
      .gout(gout),
      .pout(pout),
      .Cin(Cin),
      .g(g),
      .p(p)
   );

   overflow ov(
      .Cout(Cout),
      .V(V),
      .g(gout),
      .p(pout),
      .c31(c[31]),
      .Cin(Cin)
   );   
   
   //Zero bit 
   always @ (d) begin 
      if (d == 32'h00000000) begin
          Z = 1'b1;
      end
      else begin 
        Z = 1'b0;
      end 
   end
  
endmodule


module alu_cell (d, g, p, a, b, c, S);
   output d, g, p;
   input a, b, c;
   input [2:0] S;      
   reg g,p,d,cint,bint;
     
   always @(a,b,c,S,p,g) begin 
     bint = S[0] ^ b;
     g = a & bint;
     p = a ^ bint;
     cint = S[1] & c;
    
      if(S[2]==0)
         begin
            d = p ^ cint;
         end
         
       else if(S[2]==1)
          begin
             if((S[1]==0) & (S[0]==0)) begin
                d = a | b;
                end
             else if ((S[1]==0) & (S[0]==1)) begin
                d = ~(a | b); // nor
                end
             else if ((S[1]==1) & (S[0]==0)) begin
                d = a & b; // and 
                end   
             else
                d = 0; // undefined, but needs an output, so using 0 
                end
       end             
endmodule


module overflow (Cout, V, g, p, c31, Cin);
   output Cout, V;
   input g, p, c31, Cin;
   
   assign Cout = g|(p&Cin);
   assign V = Cout^c31;   
endmodule


module lac(c, gout, pout, Cin, g, p);

   output [1:0] c;
   output gout;
   output pout;
   input Cin;
   input [1:0] g;
   input [1:0] p;

   assign c[0] = Cin;
   assign c[1] = g[0] | ( p[0] & Cin );
   assign gout = g[1] | ( p[1] & g[0] );
   assign pout = p[1] & p[0];
	
endmodule


module lac2 (c, gout, pout, Cin, g, p);
   output [3:0] c;
   output gout, pout;
   input Cin;
   input [3:0] g, p;
   
   wire [1:0] cint, gint, pint;
   
   lac leaf0(
      .c(c[1:0]),
      .gout(gint[0]),
      .pout(pint[0]),
      .Cin(cint[0]),
      .g(g[1:0]),
      .p(p[1:0])
   );
   
   lac leaf1(
      .c(c[3:2]),
      .gout(gint[1]),
      .pout(pint[1]),
      .Cin(cint[1]),
      .g(g[3:2]),
      .p(p[3:2])
   );
   
   lac root(
      .c(cint),
      .gout(gout),
      .pout(pout),
      .Cin(Cin),
      .g(gint),
      .p(pint)
   );
endmodule   


module lac3 (c, gout, pout, Cin, g, p);
   output [7:0] c;
   output gout, pout;
   input Cin;
   input [7:0] g, p;
   
   wire [1:0] cint, gint, pint;
   
   lac2 leaf0(
      .c(c[3:0]),
      .gout(gint[0]),
      .pout(pint[0]),
      .Cin(cint[0]),
      .g(g[3:0]),
      .p(p[3:0])
   );
   
   lac2 leaf1(
      .c(c[7:4]),
      .gout(gint[1]),
      .pout(pint[1]),
      .Cin(cint[1]),
      .g(g[7:4]),
      .p(p[7:4])
   );
   
   lac root(
      .c(cint),
      .gout(gout),
      .pout(pout),
      .Cin(Cin),
      .g(gint),
      .p(pint)
   );
endmodule
      

module lac4 (c, gout, pout, Cin, g, p);
   output [15:0] c;
   output gout, pout;
   input Cin;
   input [15:0] g, p;
   
   wire [1:0] cint, gint, pint;
   
   lac3 leaf0( // First half is sent in leaf 0 
        .c(c[7:0]),
         .gout(gint[0]),
         .pout(pint[0]),
         .Cin(cint[0]),
         .g(g[7:0]),
         .p(p[7:0])
   );
   
   lac3 leaf1( // Second half is send in leaf 1 
         .c(c[15:8]),
         .gout(gint[1]),
         .pout(pint[1]),
         .Cin(cint[1]),
         .g(g[15:8]),
         .p(p[15:8])
   );
   
   lac root( // Same root as in other lacs 
      .c(cint),
      .gout(gout),
      .pout(pout),
      .Cin(Cin),
      .g(gint),
      .p(pint)
   );
endmodule
      

module lac5 (c, gout, pout, Cin, g, p);
   output [31:0] c;
   output gout, pout;
   input Cin;
   input [31:0] g, p;
   
   wire [1:0] cint, gint, pint;
   
   lac4 leaf0( // First half in leaf 0 
    .c(c[15:0]),
         .gout(gint[0]),
         .pout(pint[0]),
         .Cin(cint[0]),
         .g(g[15:0]),
         .p(p[15:0])
   );
   
   lac4 leaf1( // second half in leaf 1 
         .c(c[31:16]),
         .gout(gint[1]),
         .pout(pint[1]),
         .Cin(cint[1]),
         .g(g[31:16]),
         .p(p[31:16])
   );
   
   lac root( // Same root as in other lacs 
      .c(cint),
      .gout(gout),
      .pout(pout),
      .Cin(Cin),
      .g(gint),
      .p(pint)
   );
endmodule
